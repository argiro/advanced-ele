//-----------------------------------------------------------------------------------------------------//                               University of Torino - Department of Physics//                                   via Giuria 1 10125, Torino, Italy//-----------------------------------------------------------------------------------------------------// [Filename]       BTN_debouncer.v// [Project]        Advanced Electronics Laboratory course// [Author]         Luca Pacher - pacher@to.infn.it// [Language]       Verilog 1995 [IEEE Std. 1364-1995]// [Created]        Apr 16, 2016// [Modified]       Apr 16, 2016// [Description]    Push-button debouncer// [Notes]          -// [Version]        1.0// [Revisions]      16.04.2016 - Created//-----------------------------------------------------------------------------------------------------`timescale 1ns / 100psmodule BTN_debouncer(   input   btn,             // input pulse affected by mechanical chattering, asynchronous to clock   input   clk,      output  LE_tick,         // leading-edge and falling-edge single-pulse ticks   output  FE_tick,   output  reg pulse        // debounced output pulse      ) ;         // synchronize the input pulse with a couple of DFFs      reg btn_synch_q0, btn_synch_q1 ;      always @(posedge clk) begin      btn_synch_q0 <= btn ;      btn_synch_q1 <= btn_synch_q0 ;   end            // use a 16-bit counter to debounce the pulse      reg [15:0] btn_count ;      wire    btn_idle ;   assign  btn_idle = ( pulse == btn_synch_q1 ) ? 1'b1 : 1'b0 ;      wire   btn_count_max ;   assign btn_count_max = & btn_count ;  // carry, max. count reached      always @(posedge clk) begin         if( btn_idle )         btn_count <= 16'b0 ;      // synchronous reset !         else begin         btn_count <= btn_count + 1 ;               // output register         //if( btn_count_max )         if( btn_count == 16'hffff )            //pulse <= ~ pulse ;            pulse <= pulse ;      end // else   end // always      // assign LE/FE single-pulse ticks      assign LE_tick = (~btn_idle) & btn_count_max & (~pulse) ;   assign FE_tick = (~btn_idle) & btn_count_max & pulse ;endmodule